module testbench_pla();
    logic clk;
    logic [11:0] a;
    logic [26:0] y, expected;
    logic [38:0] vectors[27:0], currentvec;
    logic [4:0] vectornum, errors;

    // device under test
    controller_pla_Cell dut(a[0], a[1], a[10], a[11], a[2], a[3], a[4], a[5],
      a[6], a[7], a[8], a[9], y[0], y[1], y[10], y[11], y[12], y[13], 
      y[14], y[15], y[16], y[17], y[18], y[19], y[2], y[20], y[21], 
      y[22], y[23], y[24], y[25], y[26], y[3], y[4], y[5], y[6], 
      y[7], y[8], y[9]);

    // read test file and initialize test
    initial begin
        $readmemb("pla-vectors.txt", vectors);
        vectornum = 0; errors = 0;
    end
    // generate clock
    always begin
        clk = 1; #10; clk = 0; #10;
    end
    // apply test
    always @(posedge clk) begin
        currentvec = vectors[vectornum];
        a = currentvec[38:27];
        if (currentvec[0] === 1'bx) begin
            $display("Completed %d tests with %d errors.", 
                        vectornum, errors);
            $stop;
        end
    end
    // check errors
    always @(negedge clk) begin
      expected = currentvec[26:0];
        if (y !== expected) begin
            $display("       output mismatches as %h (%h expected)", 
                        y, expected);
            errors = errors + 1;
        end
        vectornum = vectornum + 1;
    end
endmodule /* testbench */

/* Verilog for cell 'controller_pla_Cell{sch}' from library 'controller_pla' */
/* Created on ÐÇÆÚÈÕ ÈýÔÂ 04, 2007 21:40:06 */
/* Last revised on ÐÇÆÚÒ» Ê®Ò»ÔÂ 17, 2014 16:41:30 */
/* Written on ÐÇÆÚÒ» Ê®Ò»ÔÂ 17, 2014 16:46:19 by Electric VLSI Design System, version 8.06 */

module controller_pla_Cell(in, in_1, in_10, in_11, in_2, in_3, in_4, in_5, 
      in_6, in_7, in_8, in_9, out, out_1, out_10, out_11, out_12, out_13, 
      out_14, out_15, out_16, out_17, out_18, out_19, out_2, out_20, out_21, 
      out_22, out_23, out_24, out_25, out_26, out_3, out_4, out_5, out_6, 
      out_7, out_8, out_9);
  input [0:0] in;
  input [1:1] in_1;
  input [10:10] in_10;
  input [11:11] in_11;
  input [2:2] in_2;
  input [3:3] in_3;
  input [4:4] in_4;
  input [5:5] in_5;
  input [6:6] in_6;
  input [7:7] in_7;
  input [8:8] in_8;
  input [9:9] in_9;
  output [0:0] out;
  output [1:1] out_1;
  output [10:10] out_10;
  output [11:11] out_11;
  output [12:12] out_12;
  output [13:13] out_13;
  output [14:14] out_14;
  output [15:15] out_15;
  output [16:16] out_16;
  output [17:17] out_17;
  output [18:18] out_18;
  output [19:19] out_19;
  output [2:2] out_2;
  output [20:20] out_20;
  output [21:21] out_21;
  output [22:22] out_22;
  output [23:23] out_23;
  output [24:24] out_24;
  output [25:25] out_25;
  output [26:26] out_26;
  output [3:3] out_3;
  output [4:4] out_4;
  output [5:5] out_5;
  output [6:6] out_6;
  output [7:7] out_7;
  output [8:8] out_8;
  output [9:9] out_9;

  supply1 vdd;
  supply0 gnd;
  wire net_0, net_1143, net_1145, net_1147, net_1149, net_1159, net_1162;
  wire net_1165, net_1168, net_1171, net_1180, net_1194, net_1196, net_1198;
  wire net_1200, net_1203, net_1207, net_1209, net_1215, net_1217, net_1228;
  wire net_1234, net_1240, net_1250, net_1263, net_1276, net_1283, net_14;
  wire net_1673, net_21, net_28, net_300, net_311, net_335, net_346, net_35;
  wire net_370, net_381, net_405, net_418, net_42, net_447, net_458, net_49;
  wire net_506, net_529, net_56, net_583, net_606, net_63, net_660, net_683;
  wire net_7, net_70, net_737, net_750, net_77, net_779, net_790, net_818;
  wire net_831, net_857, net_870, net_899, net_910, net_938, net_951;

  tranif1 nmos_3(gnd, net_0, in_11[11]);
  tranif1 nmos_10(gnd, net_7, in_10[10]);
  tranif1 nmos_17(gnd, net_14, in_9[9]);
  tranif1 nmos_24(gnd, net_21, in_8[8]);
  tranif1 nmos_31(gnd, net_28, in_7[7]);
  tranif1 nmos_38(gnd, net_35, in_6[6]);
  tranif1 nmos_45(gnd, net_42, in_5[5]);
  tranif1 nmos_52(gnd, net_49, in_4[4]);
  tranif1 nmos_59(gnd, net_56, in_3[3]);
  tranif1 nmos_66(gnd, net_63, in_2[2]);
  tranif1 nmos_73(gnd, net_70, in_1[1]);
  tranif1 nmos_80(gnd, net_77, in[0]);
  tranif1 nmos_86(net_300, gnd, in_5[5]);
  tranif1 nmos_87(net_300, gnd, net_49);
  tranif1 nmos_88(net_300, gnd, net_56);
  tranif1 nmos_89(net_300, gnd, in_2[2]);
  tranif1 nmos_90(net_300, gnd, in_1[1]);
  tranif1 nmos_91(gnd, net_311, in_5[5]);
  tranif1 nmos_92(gnd, net_311, net_49);
  tranif1 nmos_93(gnd, net_311, in_3[3]);
  tranif1 nmos_94(gnd, net_311, net_63);
  tranif1 nmos_95(gnd, net_311, net_70);
  tranif1 nmos_96(net_335, gnd, in_5[5]);
  tranif1 nmos_97(net_335, gnd, net_49);
  tranif1 nmos_98(net_335, gnd, in_3[3]);
  tranif1 nmos_99(net_335, gnd, net_63);
  tranif1 nmos_100(net_335, gnd, in_1[1]);
  tranif1 nmos_101(gnd, net_346, in_5[5]);
  tranif1 nmos_102(gnd, net_346, net_49);
  tranif1 nmos_103(gnd, net_346, in_3[3]);
  tranif1 nmos_104(gnd, net_346, in_2[2]);
  tranif1 nmos_105(gnd, net_346, net_70);
  tranif1 nmos_106(net_370, gnd, in_5[5]);
  tranif1 nmos_107(net_370, gnd, net_49);
  tranif1 nmos_108(net_370, gnd, in_3[3]);
  tranif1 nmos_109(net_370, gnd, in_2[2]);
  tranif1 nmos_110(net_370, gnd, in_1[1]);
  tranif1 nmos_111(gnd, net_381, in_5[5]);
  tranif1 nmos_112(gnd, net_381, in_4[4]);
  tranif1 nmos_113(gnd, net_381, net_56);
  tranif1 nmos_114(gnd, net_381, net_63);
  tranif1 nmos_115(gnd, net_381, net_70);
  tranif1 nmos_116(net_405, gnd, net_42);
  tranif1 nmos_117(net_405, gnd, in_4[4]);
  tranif1 nmos_118(net_405, gnd, net_56);
  tranif1 nmos_119(net_405, gnd, net_63);
  tranif1 nmos_120(net_405, gnd, in_1[1]);
  tranif1 nmos_121(net_405, gnd, net_77);
  tranif1 nmos_122(gnd, net_418, net_42);
  tranif1 nmos_123(gnd, net_418, in_4[4]);
  tranif1 nmos_124(gnd, net_418, net_56);
  tranif1 nmos_125(gnd, net_418, net_63);
  tranif1 nmos_126(gnd, net_418, in_1[1]);
  tranif1 nmos_127(gnd, net_418, in[0]);
  tranif1 nmos_128(net_447, gnd, in_5[5]);
  tranif1 nmos_129(net_447, gnd, in_4[4]);
  tranif1 nmos_130(net_447, gnd, net_56);
  tranif1 nmos_131(net_447, gnd, net_63);
  tranif1 nmos_132(net_447, gnd, in_1[1]);
  tranif1 nmos_133(gnd, net_458, net_0);
  tranif1 nmos_134(gnd, net_458, in_10[10]);
  tranif1 nmos_135(gnd, net_458, net_14);
  tranif1 nmos_136(gnd, net_458, in_8[8]);
  tranif1 nmos_137(gnd, net_458, in_7[7]);
  tranif1 nmos_138(gnd, net_458, in_6[6]);
  tranif1 nmos_139(gnd, net_458, in_5[5]);
  tranif1 nmos_140(gnd, net_458, in_4[4]);
  tranif1 nmos_141(gnd, net_458, net_56);
  tranif1 nmos_142(gnd, net_458, in_2[2]);
  tranif1 nmos_143(gnd, net_458, net_70);
  tranif1 nmos_144(net_506, gnd, net_0);
  tranif1 nmos_145(net_506, gnd, in_10[10]);
  tranif1 nmos_146(net_506, gnd, in_9[9]);
  tranif1 nmos_147(net_506, gnd, in_8[8]);
  tranif1 nmos_148(net_506, gnd, in_7[7]);
  tranif1 nmos_149(net_506, gnd, in_6[6]);
  tranif1 nmos_150(net_506, gnd, in_5[5]);
  tranif1 nmos_151(net_506, gnd, in_4[4]);
  tranif1 nmos_152(net_506, gnd, net_56);
  tranif1 nmos_153(net_506, gnd, in_2[2]);
  tranif1 nmos_154(net_506, gnd, net_70);
  tranif1 nmos_155(gnd, net_529, in_11[11]);
  tranif1 nmos_156(gnd, net_529, in_10[10]);
  tranif1 nmos_157(gnd, net_529, in_9[9]);
  tranif1 nmos_158(gnd, net_529, in_8[8]);
  tranif1 nmos_159(gnd, net_529, net_28);
  tranif1 nmos_160(gnd, net_529, in_6[6]);
  tranif1 nmos_161(gnd, net_529, in_5[5]);
  tranif1 nmos_162(gnd, net_529, in_4[4]);
  tranif1 nmos_163(gnd, net_529, net_56);
  tranif1 nmos_164(gnd, net_529, in_2[2]);
  tranif1 nmos_165(gnd, net_529, in_1[1]);
  tranif1 nmos_166(net_583, gnd, in_11[11]);
  tranif1 nmos_167(net_583, gnd, in_10[10]);
  tranif1 nmos_168(net_583, gnd, in_9[9]);
  tranif1 nmos_169(net_583, gnd, net_21);
  tranif1 nmos_170(net_583, gnd, in_7[7]);
  tranif1 nmos_171(net_583, gnd, in_6[6]);
  tranif1 nmos_172(net_583, gnd, in_5[5]);
  tranif1 nmos_173(net_583, gnd, in_4[4]);
  tranif1 nmos_174(net_583, gnd, net_56);
  tranif1 nmos_175(net_583, gnd, in_2[2]);
  tranif1 nmos_176(net_583, gnd, in_1[1]);
  tranif1 nmos_177(gnd, net_606, in_11[11]);
  tranif1 nmos_178(gnd, net_606, in_10[10]);
  tranif1 nmos_179(gnd, net_606, in_9[9]);
  tranif1 nmos_180(gnd, net_606, in_8[8]);
  tranif1 nmos_181(gnd, net_606, in_7[7]);
  tranif1 nmos_182(gnd, net_606, in_6[6]);
  tranif1 nmos_183(gnd, net_606, in_5[5]);
  tranif1 nmos_184(gnd, net_606, in_4[4]);
  tranif1 nmos_185(gnd, net_606, net_56);
  tranif1 nmos_186(gnd, net_606, in_2[2]);
  tranif1 nmos_187(gnd, net_606, in_1[1]);
  tranif1 nmos_188(net_660, gnd, net_0);
  tranif1 nmos_189(net_660, gnd, in_10[10]);
  tranif1 nmos_190(net_660, gnd, net_14);
  tranif1 nmos_191(net_660, gnd, in_8[8]);
  tranif1 nmos_192(net_660, gnd, in_7[7]);
  tranif1 nmos_193(net_660, gnd, in_6[6]);
  tranif1 nmos_194(net_660, gnd, in_5[5]);
  tranif1 nmos_195(net_660, gnd, in_4[4]);
  tranif1 nmos_196(net_660, gnd, net_56);
  tranif1 nmos_197(net_660, gnd, in_2[2]);
  tranif1 nmos_198(net_660, gnd, in_1[1]);
  tranif1 nmos_199(gnd, net_683, net_0);
  tranif1 nmos_200(gnd, net_683, in_10[10]);
  tranif1 nmos_201(gnd, net_683, in_9[9]);
  tranif1 nmos_202(gnd, net_683, in_8[8]);
  tranif1 nmos_203(gnd, net_683, in_7[7]);
  tranif1 nmos_204(gnd, net_683, in_6[6]);
  tranif1 nmos_205(gnd, net_683, in_5[5]);
  tranif1 nmos_206(gnd, net_683, in_4[4]);
  tranif1 nmos_207(gnd, net_683, net_56);
  tranif1 nmos_208(gnd, net_683, in_2[2]);
  tranif1 nmos_209(gnd, net_683, in_1[1]);
  tranif1 nmos_210(net_737, gnd, net_42);
  tranif1 nmos_211(net_737, gnd, in_4[4]);
  tranif1 nmos_212(net_737, gnd, in_3[3]);
  tranif1 nmos_213(net_737, gnd, net_63);
  tranif1 nmos_214(net_737, gnd, net_70);
  tranif1 nmos_215(net_737, gnd, net_77);
  tranif1 nmos_216(gnd, net_750, net_42);
  tranif1 nmos_217(gnd, net_750, in_4[4]);
  tranif1 nmos_218(gnd, net_750, in_3[3]);
  tranif1 nmos_219(gnd, net_750, net_63);
  tranif1 nmos_220(gnd, net_750, net_70);
  tranif1 nmos_221(gnd, net_750, in[0]);
  tranif1 nmos_222(net_779, gnd, in_5[5]);
  tranif1 nmos_223(net_779, gnd, in_4[4]);
  tranif1 nmos_224(net_779, gnd, in_3[3]);
  tranif1 nmos_225(net_779, gnd, net_63);
  tranif1 nmos_226(net_779, gnd, net_70);
  tranif1 nmos_227(gnd, net_790, net_42);
  tranif1 nmos_228(gnd, net_790, in_4[4]);
  tranif1 nmos_229(gnd, net_790, in_3[3]);
  tranif1 nmos_230(gnd, net_790, net_63);
  tranif1 nmos_231(gnd, net_790, in_1[1]);
  tranif1 nmos_232(gnd, net_790, net_77);
  tranif1 nmos_233(net_818, gnd, net_42);
  tranif1 nmos_234(net_818, gnd, in_4[4]);
  tranif1 nmos_235(net_818, gnd, in_3[3]);
  tranif1 nmos_236(net_818, gnd, net_63);
  tranif1 nmos_237(net_818, gnd, in_1[1]);
  tranif1 nmos_238(net_818, gnd, in[0]);
  tranif1 nmos_239(gnd, net_831, in_5[5]);
  tranif1 nmos_240(gnd, net_831, in_4[4]);
  tranif1 nmos_241(gnd, net_831, in_3[3]);
  tranif1 nmos_242(gnd, net_831, net_63);
  tranif1 nmos_243(gnd, net_831, in_1[1]);
  tranif1 nmos_244(net_857, gnd, net_42);
  tranif1 nmos_245(net_857, gnd, in_4[4]);
  tranif1 nmos_246(net_857, gnd, in_3[3]);
  tranif1 nmos_247(net_857, gnd, in_2[2]);
  tranif1 nmos_248(net_857, gnd, net_70);
  tranif1 nmos_249(net_857, gnd, net_77);
  tranif1 nmos_250(gnd, net_870, net_42);
  tranif1 nmos_251(gnd, net_870, in_4[4]);
  tranif1 nmos_252(gnd, net_870, in_3[3]);
  tranif1 nmos_253(gnd, net_870, in_2[2]);
  tranif1 nmos_254(gnd, net_870, net_70);
  tranif1 nmos_255(gnd, net_870, in[0]);
  tranif1 nmos_256(net_899, gnd, in_5[5]);
  tranif1 nmos_257(net_899, gnd, in_4[4]);
  tranif1 nmos_258(net_899, gnd, in_3[3]);
  tranif1 nmos_259(net_899, gnd, in_2[2]);
  tranif1 nmos_260(net_899, gnd, net_70);
  tranif1 nmos_261(gnd, net_910, net_42);
  tranif1 nmos_262(gnd, net_910, in_4[4]);
  tranif1 nmos_263(gnd, net_910, in_3[3]);
  tranif1 nmos_264(gnd, net_910, in_2[2]);
  tranif1 nmos_265(gnd, net_910, in_1[1]);
  tranif1 nmos_266(gnd, net_910, net_77);
  tranif1 nmos_267(net_938, gnd, net_42);
  tranif1 nmos_268(net_938, gnd, in_4[4]);
  tranif1 nmos_269(net_938, gnd, in_3[3]);
  tranif1 nmos_270(net_938, gnd, in_2[2]);
  tranif1 nmos_271(net_938, gnd, in_1[1]);
  tranif1 nmos_272(net_938, gnd, in[0]);
  tranif1 nmos_273(gnd, net_951, in_5[5]);
  tranif1 nmos_274(gnd, net_951, in_4[4]);
  tranif1 nmos_275(gnd, net_951, in_3[3]);
  tranif1 nmos_276(gnd, net_951, in_2[2]);
  tranif1 nmos_277(gnd, net_951, in_1[1]);
  tranif1 nmos_646(gnd, net_1149, net_300);
  tranif1 nmos_647(gnd, net_1194, net_300);
  tranif1 nmos_648(gnd, net_1145, net_311);
  tranif1 nmos_649(gnd, net_1147, net_311);
  tranif1 nmos_650(gnd, net_1196, net_311);
  tranif1 nmos_651(gnd, net_1209, net_311);
  tranif1 nmos_652(gnd, net_1198, net_335);
  tranif1 nmos_653(gnd, net_1200, net_335);
  tranif1 nmos_654(gnd, net_1143, net_346);
  tranif1 nmos_655(gnd, net_1209, net_346);
  tranif1 nmos_656(gnd, net_1234, net_346);
  tranif1 nmos_657(gnd, net_1250, net_346);
  tranif1 nmos_658(gnd, net_1203, net_370);
  tranif1 nmos_659(gnd, net_1215, net_370);
  tranif1 nmos_660(gnd, net_1276, net_370);
  tranif1 nmos_661(gnd, net_1200, net_381);
  tranif1 nmos_662(gnd, net_1207, net_381);
  tranif1 nmos_663(gnd, net_1203, net_405);
  tranif1 nmos_664(gnd, net_1217, net_405);
  tranif1 nmos_665(gnd, net_1240, net_405);
  tranif1 nmos_666(gnd, net_1250, net_405);
  tranif1 nmos_667(gnd, net_1263, net_405);
  tranif1 nmos_668(gnd, net_1283, net_405);
  tranif1 nmos_669(gnd, net_1203, net_418);
  tranif1 nmos_670(gnd, net_1217, net_418);
  tranif1 nmos_671(gnd, net_1240, net_418);
  tranif1 nmos_672(gnd, net_1250, net_418);
  tranif1 nmos_673(gnd, net_1263, net_418);
  tranif1 nmos_674(gnd, net_1276, net_418);
  tranif1 nmos_675(gnd, net_1171, net_447);
  tranif1 nmos_676(gnd, net_1209, net_447);
  tranif1 nmos_677(gnd, net_1228, net_447);
  tranif1 nmos_678(gnd, net_1240, net_447);
  tranif1 nmos_679(gnd, net_1250, net_447);
  tranif1 nmos_680(gnd, net_1171, net_458);
  tranif1 nmos_681(gnd, net_1209, net_458);
  tranif1 nmos_682(gnd, net_1234, net_458);
  tranif1 nmos_683(gnd, net_1171, net_506);
  tranif1 nmos_684(gnd, net_1209, net_506);
  tranif1 nmos_685(gnd, net_1240, net_506);
  tranif1 nmos_686(gnd, net_1250, net_506);
  tranif1 nmos_687(gnd, net_1171, net_529);
  tranif1 nmos_688(gnd, net_1180, net_529);
  tranif1 nmos_689(gnd, net_1234, net_529);
  tranif1 nmos_690(gnd, net_1240, net_529);
  tranif1 nmos_691(gnd, net_1171, net_583);
  tranif1 nmos_692(gnd, net_1180, net_583);
  tranif1 nmos_693(gnd, net_1234, net_583);
  tranif1 nmos_694(gnd, net_1250, net_583);
  tranif1 nmos_695(gnd, net_1263, net_583);
  tranif1 nmos_696(gnd, net_1171, net_606);
  tranif1 nmos_697(gnd, net_1180, net_606);
  tranif1 nmos_698(gnd, net_1234, net_606);
  tranif1 nmos_699(gnd, net_1263, net_606);
  tranif1 nmos_700(gnd, net_1171, net_660);
  tranif1 nmos_701(gnd, net_1180, net_660);
  tranif1 nmos_702(gnd, net_1240, net_660);
  tranif1 nmos_703(gnd, net_1263, net_660);
  tranif1 nmos_704(gnd, net_1171, net_683);
  tranif1 nmos_705(gnd, net_1180, net_683);
  tranif1 nmos_706(gnd, net_1240, net_683);
  tranif1 nmos_707(gnd, net_1263, net_683);
  tranif1 nmos_708(gnd, net_1149, net_737);
  tranif1 nmos_709(gnd, net_1159, net_737);
  tranif1 nmos_710(gnd, net_1180, net_737);
  tranif1 nmos_711(gnd, net_1217, net_737);
  tranif1 nmos_712(gnd, net_1240, net_737);
  tranif1 nmos_713(gnd, net_1283, net_737);
  tranif1 nmos_714(gnd, net_1149, net_750);
  tranif1 nmos_715(gnd, net_1159, net_750);
  tranif1 nmos_716(gnd, net_1180, net_750);
  tranif1 nmos_717(gnd, net_1217, net_750);
  tranif1 nmos_718(gnd, net_1240, net_750);
  tranif1 nmos_719(gnd, net_1276, net_750);
  tranif1 nmos_720(gnd, net_1228, net_779);
  tranif1 nmos_721(gnd, net_1250, net_779);
  tranif1 nmos_722(gnd, net_1263, net_779);
  tranif1 nmos_723(gnd, net_1149, net_790);
  tranif1 nmos_724(gnd, net_1162, net_790);
  tranif1 nmos_725(gnd, net_1180, net_790);
  tranif1 nmos_726(gnd, net_1217, net_790);
  tranif1 nmos_727(gnd, net_1250, net_790);
  tranif1 nmos_728(gnd, net_1263, net_790);
  tranif1 nmos_729(gnd, net_1283, net_790);
  tranif1 nmos_730(gnd, net_1149, net_818);
  tranif1 nmos_731(gnd, net_1162, net_818);
  tranif1 nmos_732(gnd, net_1180, net_818);
  tranif1 nmos_733(gnd, net_1217, net_818);
  tranif1 nmos_734(gnd, net_1250, net_818);
  tranif1 nmos_735(gnd, net_1263, net_818);
  tranif1 nmos_736(gnd, net_1276, net_818);
  tranif1 nmos_737(gnd, net_1228, net_831);
  tranif1 nmos_738(gnd, net_1250, net_831);
  tranif1 nmos_739(gnd, net_1149, net_857);
  tranif1 nmos_740(gnd, net_1165, net_857);
  tranif1 nmos_741(gnd, net_1180, net_857);
  tranif1 nmos_742(gnd, net_1217, net_857);
  tranif1 nmos_743(gnd, net_1250, net_857);
  tranif1 nmos_744(gnd, net_1283, net_857);
  tranif1 nmos_745(gnd, net_1149, net_870);
  tranif1 nmos_746(gnd, net_1165, net_870);
  tranif1 nmos_747(gnd, net_1180, net_870);
  tranif1 nmos_748(gnd, net_1217, net_870);
  tranif1 nmos_749(gnd, net_1250, net_870);
  tranif1 nmos_750(gnd, net_1276, net_870);
  tranif1 nmos_751(gnd, net_1228, net_899);
  tranif1 nmos_752(gnd, net_1263, net_899);
  tranif1 nmos_753(gnd, net_1149, net_910);
  tranif1 nmos_754(gnd, net_1168, net_910);
  tranif1 nmos_755(gnd, net_1180, net_910);
  tranif1 nmos_756(gnd, net_1217, net_910);
  tranif1 nmos_757(gnd, net_1263, net_910);
  tranif1 nmos_758(gnd, net_1283, net_910);
  tranif1 nmos_759(gnd, net_1149, net_938);
  tranif1 nmos_760(gnd, net_1168, net_938);
  tranif1 nmos_761(gnd, net_1180, net_938);
  tranif1 nmos_762(gnd, net_1217, net_938);
  tranif1 nmos_763(gnd, net_1263, net_938);
  tranif1 nmos_764(gnd, net_1276, net_938);
  tranif1 nmos_765(gnd, net_1228, net_951);
  tranif1 nmos_878(gnd, out_26[26], net_1143);
  tranif1 nmos_886(gnd, out_25[25], net_1145);
  tranif1 nmos_894(gnd, out_24[24], net_1147);
  tranif1 nmos_902(gnd, out_23[23], net_1149);
  tranif1 nmos_910(gnd, out_22[22], net_1159);
  tranif1 nmos_918(gnd, out_21[21], net_1162);
  tranif1 nmos_926(gnd, out_20[20], net_1165);
  tranif1 nmos_934(gnd, out_19[19], net_1168);
  tranif1 nmos_942(gnd, out_18[18], net_1171);
  tranif1 nmos_950(gnd, out_17[17], net_1180);
  tranif1 nmos_958(gnd, out_16[16], net_1194);
  tranif1 nmos_966(gnd, out_15[15], net_1196);
  tranif1 nmos_974(gnd, out_14[14], net_1198);
  tranif1 nmos_982(gnd, out_13[13], net_1200);
  tranif1 nmos_990(gnd, out_12[12], net_1203);
  tranif1 nmos_998(gnd, out_11[11], net_1207);
  tranif1 nmos_1006(gnd, out_10[10], net_1209);
  tranif1 nmos_1014(gnd, out_9[9], net_1215);
  tranif1 nmos_1022(gnd, out_8[8], net_1217);
  tranif1 nmos_1030(gnd, out_7[7], net_1228);
  tranif1 nmos_1038(gnd, out_6[6], net_1234);
  tranif1 nmos_1046(gnd, out_5[5], net_1240);
  tranif1 nmos_1054(gnd, out_4[4], net_1250);
  tranif1 nmos_1062(gnd, out_3[3], net_1263);
  tranif1 nmos_1070(gnd, out_2[2], net_1276);
  tranif1 nmos_1078(gnd, out_1[1], net_1283);
  tranif1 nmos_1086(gnd, out[0], net_1673);
  tranif0 pmos_4(net_0, vdd, in_11[11]);
  tranif0 pmos_11(net_7, vdd, in_10[10]);
  tranif0 pmos_18(net_14, vdd, in_9[9]);
  tranif0 pmos_25(net_21, vdd, in_8[8]);
  tranif0 pmos_32(net_28, vdd, in_7[7]);
  tranif0 pmos_39(net_35, vdd, in_6[6]);
  tranif0 pmos_46(net_42, vdd, in_5[5]);
  tranif0 pmos_53(net_49, vdd, in_4[4]);
  tranif0 pmos_60(net_56, vdd, in_3[3]);
  tranif0 pmos_67(net_63, vdd, in_2[2]);
  tranif0 pmos_74(net_70, vdd, in_1[1]);
  tranif0 pmos_81(net_77, vdd, in[0]);
  tranif0 pmos_879(out_26[26], vdd, net_1143);
  tranif0 pmos_887(out_25[25], vdd, net_1145);
  tranif0 pmos_895(out_24[24], vdd, net_1147);
  tranif0 pmos_903(out_23[23], vdd, net_1149);
  tranif0 pmos_911(out_22[22], vdd, net_1159);
  tranif0 pmos_919(out_21[21], vdd, net_1162);
  tranif0 pmos_927(out_20[20], vdd, net_1165);
  tranif0 pmos_935(out_19[19], vdd, net_1168);
  tranif0 pmos_943(out_18[18], vdd, net_1171);
  tranif0 pmos_951(out_17[17], vdd, net_1180);
  tranif0 pmos_959(out_16[16], vdd, net_1194);
  tranif0 pmos_967(out_15[15], vdd, net_1196);
  tranif0 pmos_975(out_14[14], vdd, net_1198);
  tranif0 pmos_983(out_13[13], vdd, net_1200);
  tranif0 pmos_991(out_12[12], vdd, net_1203);
  tranif0 pmos_999(out_11[11], vdd, net_1207);
  tranif0 pmos_1007(out_10[10], vdd, net_1209);
  tranif0 pmos_1015(out_9[9], vdd, net_1215);
  tranif0 pmos_1023(out_8[8], vdd, net_1217);
  tranif0 pmos_1031(out_7[7], vdd, net_1228);
  tranif0 pmos_1039(out_6[6], vdd, net_1234);
  tranif0 pmos_1047(out_5[5], vdd, net_1240);
  tranif0 pmos_1055(out_4[4], vdd, net_1250);
  tranif0 pmos_1063(out_3[3], vdd, net_1263);
  tranif0 pmos_1071(out_2[2], vdd, net_1276);
  tranif0 pmos_1079(out_1[1], vdd, net_1283);
  tranif0 pmos_1087(out[0], vdd, net_1673);
  rtranif0 pmos_1092(net_1143, vdd, gnd);
  rtranif0 pmos_1094(net_1145, vdd, gnd);
  rtranif0 pmos_1096(net_1147, vdd, gnd);
  rtranif0 pmos_1098(net_1149, vdd, gnd);
  rtranif0 pmos_1100(net_1159, vdd, gnd);
  rtranif0 pmos_1102(net_1162, vdd, gnd);
  rtranif0 pmos_1104(net_1165, vdd, gnd);
  rtranif0 pmos_1106(net_1168, vdd, gnd);
  rtranif0 pmos_1108(net_1171, vdd, gnd);
  rtranif0 pmos_1110(net_1180, vdd, gnd);
  rtranif0 pmos_1112(net_1194, vdd, gnd);
  rtranif0 pmos_1114(net_1196, vdd, gnd);
  rtranif0 pmos_1116(net_1198, vdd, gnd);
  rtranif0 pmos_1118(net_1200, vdd, gnd);
  rtranif0 pmos_1120(net_1203, vdd, gnd);
  rtranif0 pmos_1122(net_1207, vdd, gnd);
  rtranif0 pmos_1124(net_1209, vdd, gnd);
  rtranif0 pmos_1126(net_1215, vdd, gnd);
  rtranif0 pmos_1128(net_1217, vdd, gnd);
  rtranif0 pmos_1130(net_1228, vdd, gnd);
  rtranif0 pmos_1132(net_1234, vdd, gnd);
  rtranif0 pmos_1134(net_1240, vdd, gnd);
  rtranif0 pmos_1136(net_1250, vdd, gnd);
  rtranif0 pmos_1138(net_1263, vdd, gnd);
  rtranif0 pmos_1140(net_1276, vdd, gnd);
  rtranif0 pmos_1142(net_1283, vdd, gnd);
  rtranif0 pmos_1144(net_1673, vdd, gnd);
  rtranif0 pmos_1148(vdd, net_951, gnd);
  rtranif0 pmos_1150(vdd, net_938, gnd);
  rtranif0 pmos_1152(vdd, net_910, gnd);
  rtranif0 pmos_1154(vdd, net_899, gnd);
  rtranif0 pmos_1156(vdd, net_870, gnd);
  rtranif0 pmos_1158(vdd, net_857, gnd);
  rtranif0 pmos_1160(vdd, net_831, gnd);
  rtranif0 pmos_1162(vdd, net_818, gnd);
  rtranif0 pmos_1164(vdd, net_790, gnd);
  rtranif0 pmos_1166(vdd, net_779, gnd);
  rtranif0 pmos_1168(vdd, net_750, gnd);
  rtranif0 pmos_1170(vdd, net_737, gnd);
  rtranif0 pmos_1172(vdd, net_683, gnd);
  rtranif0 pmos_1174(vdd, net_660, gnd);
  rtranif0 pmos_1176(vdd, net_606, gnd);
  rtranif0 pmos_1178(vdd, net_583, gnd);
  rtranif0 pmos_1180(vdd, net_529, gnd);
  rtranif0 pmos_1182(vdd, net_506, gnd);
  rtranif0 pmos_1184(vdd, net_458, gnd);
  rtranif0 pmos_1186(vdd, net_447, gnd);
  rtranif0 pmos_1188(vdd, net_418, gnd);
  rtranif0 pmos_1190(vdd, net_405, gnd);
  rtranif0 pmos_1192(vdd, net_381, gnd);
  rtranif0 pmos_1194(vdd, net_370, gnd);
  rtranif0 pmos_1196(vdd, net_346, gnd);
  rtranif0 pmos_1198(vdd, net_335, gnd);
  rtranif0 pmos_1200(vdd, net_311, gnd);
  rtranif0 pmos_1202(vdd, net_300, gnd);
endmodule   /* controller_pla_Cell */
