*** SPICE deck for cell and2_1x{sch} from library muddlib07
*** Created on ������ һ�� 25, 2007 11:45:29
*** Last revised on ����һ ���� 12, 2007 05:28:50
*** Written on ������ ʮһ�� 27, 2014 23:29:29 by Electric VLSI Design System, 
*version 8.06
*** Layout tech: mocmos, foundry MOSIS
*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF
.MODEL N NMOS LEVEL=2 LD=0.3943U TOX=502E-10
+NSUB=1.22416E+16 VTO=0.756 KP=4.224E-05 GAMMA=0.9241
+PHI=0.6 UO=623.661 UEXP=8.328627E-02 UCRIT=54015.0
+DELTA=5.218409E-03 VMAX=50072.2 XJ=0.4U LAMBDA=2.975321E-02
+NFS=4.909947E+12 NEFF=1.001E-02 NSS=0.0 TPG=1.0
+RSH=20.37 CGDO=3.1E-10 CGSO=3.1E-10
+CJ=3.205E-04 MJ=0.4579 CJSW=4.62E-10 MJSW=0.2955 PB=0.7
.MODEL P PMOS LEVEL=2 LD=0.2875U TOX=502E-10
+NSUB=1.715148E+15 VTO=-0.7045 KP=1.686E-05 GAMMA=0.3459
+PHI=0.6 UO=248.933 UEXP=1.02652 UCRIT=182055.0
+DELTA=1.0E-06 VMAX=100000.0 XJ=0.4U LAMBDA=1.25919E-02
+NFS=1.0E+12 NEFF=1.001E-02 NSS=0.0 TPG=-1.0
+RSH=79.10 CGDO=2.89E-10 CGSO=2.89E-10
+CJ=1.319E-04 MJ=0.4125 CJSW=3.421E-10 MJSW=0.198 PB=0.66
.TEMP 25.0

*** TOP LEVEL CELL: muddlib07:and2_1x{sch}
Mnmos_0 net_2 b net_1 0 N L=1.2U W=3.6U
Mnmos_1 net_1 a 0 0 N L=1.2U W=3.6U
Mnmos_2 y net_2 0 0 N L=1.2U W=4.2U
Mpmos_0 vdd b net_2 vdd P L=1.2U W=3.6U
Mpmos_1 vdd a net_2 vdd P L=1.2U W=3.6U
Mpmos_2 vdd net_2 y vdd P L=1.2U W=6U

Vdd vdd 0 DC 5
*Va a 0 DC 5
Va a 0 PULSE(0 5 1u 20u 20u 480u 1m)
Vb b 0 DC 5
*Rb b 0 1k

.TRAN 1u 5m 0 1u
.PROBE

.END
